
module System2M (
	clk_cpu_clk,
	reset_reset_n);	

	input		clk_cpu_clk;
	input		reset_reset_n;
endmodule
